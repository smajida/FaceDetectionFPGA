-- megafunction wizard: %ALTSQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTSQRT 

-- ============================================================
-- File Name: altsqrt_unsign54bit_to_usign54bit.vhd
-- Megafunction Name(s):
-- 			ALTSQRT
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 14.1.0 Build 186 12/03/2014 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY altsqrt_unsign54bit_to_usign54bit IS
	PORT
	(
		radical		: IN STD_LOGIC_VECTOR (53 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
		remainder		: OUT STD_LOGIC_VECTOR (27 DOWNTO 0)
	);
END altsqrt_unsign54bit_to_usign54bit;


ARCHITECTURE SYN OF altsqrt_unsign54bit_to_usign54bit IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (26 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (27 DOWNTO 0);



	COMPONENT altsqrt
	GENERIC (
		pipeline		: NATURAL;
		q_port_width		: NATURAL;
		r_port_width		: NATURAL;
		width		: NATURAL;
		lpm_type		: STRING
	);
	PORT (
			radical	: IN STD_LOGIC_VECTOR (53 DOWNTO 0);
			q	: OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
			remainder	: OUT STD_LOGIC_VECTOR (27 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(26 DOWNTO 0);
	remainder    <= sub_wire1(27 DOWNTO 0);

	ALTSQRT_component : ALTSQRT
	GENERIC MAP (
		pipeline => 0,
		q_port_width => 27,
		r_port_width => 28,
		width => 54,
		lpm_type => "ALTSQRT"
	)
	PORT MAP (
		radical => radical,
		q => sub_wire0,
		remainder => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "27"
-- Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "28"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "54"
-- Retrieval info: USED_PORT: q 0 0 27 0 OUTPUT NODEFVAL "q[26..0]"
-- Retrieval info: USED_PORT: radical 0 0 54 0 INPUT NODEFVAL "radical[53..0]"
-- Retrieval info: USED_PORT: remainder 0 0 28 0 OUTPUT NODEFVAL "remainder[27..0]"
-- Retrieval info: CONNECT: @radical 0 0 54 0 radical 0 0 54 0
-- Retrieval info: CONNECT: q 0 0 27 0 @q 0 0 27 0
-- Retrieval info: CONNECT: remainder 0 0 28 0 @remainder 0 0 28 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_unsign54bit_to_usign54bit.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_unsign54bit_to_usign54bit.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_unsign54bit_to_usign54bit.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_unsign54bit_to_usign54bit.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_unsign54bit_to_usign54bit_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
